library IEEE;
use IEEE.std_logic_1164.all;
use ieee.numeric_std.ALL;
use work.perceptron.all;

entity fp_matrix_multiplication is
	generic(
		A_row : integer := 2;
		A_column : integer := 2;
		B_row : integer := 2;
		B_column :integer := 2;		
		i_bits : integer := 32);
	port( A : in std_logic_vector((A_row*A_column*i_bits)-1 downto 0); 
			B : in std_logic_vector((B_row*B_column*i_bits)-1 downto 0);
			c : OUT std_logic_vector((A_column*B_row*(i_bits))-1 downto 0)); --multiplication is A x B
end fp_matrix_multiplication;

architecture behavioral of fp_matrix_multiplication is

	--intermediate matrix format
	type A_matrixType is array(0 to A_row-1, 0 to A_column-1) of std_logic_vector(i_bits-1 downto 0);
	signal matA : A_matrixType;
	type B_matrixType is array(0 to B_row-1, 0 to B_column-1) of std_logic_vector(i_bits-1 downto 0);
	signal matB : B_matrixType;
	signal i, j, k: integer :=0;
	type outType is array(0 to A_column-1, 0 to B_row-1) of std_logic_vector((i_bits)-1 downto 0);
	signal matC : outType ;
	
	signal mult_temp : std_logic_vector(i_bits-1 downto 0);
	signal element : std_logic_vector((i_bits)-1 downto 0);
	signal inter : std_logic_vector((i_bits)-1 downto 0);
		
	begin
	
	inter <= (others => '0');
	
	process (A, B, matA, matB, matC)
		begin
		for i in 0 to A_row-1 loop
			for j in 0 to A_column-1 loop
				matA(i,j) <= A(((i*A_row+j+1)*i_bits)-1 downto (i*A_row+j)*i_bits);
			end loop;
		end loop;
		
		for i in 0 to B_row-1 loop
			for j in 0 to B_column-1 loop
				matB(i,j) <= B(((i*B_row+j+1)*i_bits)-1 downto (i*B_row+j)*i_bits);
			end loop;
		end loop;
	end process;		
						
	--multiplication of 2D matrix
	FA_BANK1:
	for i in 0 to A_column-1 generate --matC_row
		FA_BANK2:
		for j in 0 to B_row-1 generate --matC_column
			FA_BANK3:
			for k in 0 to B_row-1 generate --either B_row ==A_column
				M1 : multiplication_fp_general port map(matA(i,k), matB(k,j), mult_temp);
				inter <= std_logic_vector( unsigned(inter) + unsigned(mult_temp));
			end generate;
			matC(i,j) <= inter;
		end generate;
	end generate;
		
	process (A, B, matA, matB, matC)
		begin
		--return in 1D matrix
		for i in 0 to B_column-1 loop --matC_row
			for j in 0 to A_row-1 loop --matC_column
				element <= matC(i,j);
				C(((i*B_column+j+1)*(i_bits)-1) downto (i*B_column+j)*(i_bits)) <= element;
			end loop;
		end loop;
	end process;
	
end architecture;

